// lab3_qsys.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module lab3_qsys (
		input  wire       clk_clk,                                  //                               clk.clk
		output wire [3:0] digit0_external_connection_export,        //        digit0_external_connection.export
		output wire [3:0] digit1_external_connection_export,        //        digit1_external_connection.export
		output wire [3:0] digit2_external_connection_export,        //        digit2_external_connection.export
		output wire [3:0] digit3_external_connection_export,        //        digit3_external_connection.export
		output wire [3:0] digit4_external_connection_export,        //        digit4_external_connection.export
		output wire [3:0] digit5_external_connection_export,        //        digit5_external_connection.export
		inout  wire       opencores_i2c_0_export_0_scl_pad_io,      //          opencores_i2c_0_export_0.scl_pad_io
		inout  wire       opencores_i2c_0_export_0_sda_pad_io,      //                                  .sda_pad_io
		input  wire       piopushbutton_external_connection_export, // piopushbutton_external_connection.export
		input  wire       reset_reset_n                             //                             reset.reset_n
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                            // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                         // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [17:0] nios2_gen2_0_data_master_address;                             // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                          // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                               // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                           // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [17:0] nios2_gen2_0_instruction_master_address;                      // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                         // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect;  // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_chipselect -> opencores_i2c_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata;    // opencores_i2c_0:wb_dat_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest; // opencores_i2c_0:wb_ack_o -> mm_interconnect_0:opencores_i2c_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address;     // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_address -> opencores_i2c_0:wb_adr_i
	wire         mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write;       // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_write -> opencores_i2c_0:wb_we_i
	wire   [7:0] mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata;   // mm_interconnect_0:opencores_i2c_0_avalon_slave_0_writedata -> opencores_i2c_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;      // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;   // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                  // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_s1_address;                   // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                     // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                 // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                     // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_digit0_s1_chipselect;                       // mm_interconnect_0:digit0_s1_chipselect -> digit0:chipselect
	wire  [31:0] mm_interconnect_0_digit0_s1_readdata;                         // digit0:readdata -> mm_interconnect_0:digit0_s1_readdata
	wire   [2:0] mm_interconnect_0_digit0_s1_address;                          // mm_interconnect_0:digit0_s1_address -> digit0:address
	wire         mm_interconnect_0_digit0_s1_write;                            // mm_interconnect_0:digit0_s1_write -> digit0:write_n
	wire  [31:0] mm_interconnect_0_digit0_s1_writedata;                        // mm_interconnect_0:digit0_s1_writedata -> digit0:writedata
	wire         mm_interconnect_0_piopushbutton_s1_chipselect;                // mm_interconnect_0:pioPushButton_s1_chipselect -> pioPushButton:chipselect
	wire  [31:0] mm_interconnect_0_piopushbutton_s1_readdata;                  // pioPushButton:readdata -> mm_interconnect_0:pioPushButton_s1_readdata
	wire   [1:0] mm_interconnect_0_piopushbutton_s1_address;                   // mm_interconnect_0:pioPushButton_s1_address -> pioPushButton:address
	wire         mm_interconnect_0_piopushbutton_s1_write;                     // mm_interconnect_0:pioPushButton_s1_write -> pioPushButton:write_n
	wire  [31:0] mm_interconnect_0_piopushbutton_s1_writedata;                 // mm_interconnect_0:pioPushButton_s1_writedata -> pioPushButton:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                        // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                          // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                           // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                             // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                         // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_digit1_s1_chipselect;                       // mm_interconnect_0:digit1_s1_chipselect -> digit1:chipselect
	wire  [31:0] mm_interconnect_0_digit1_s1_readdata;                         // digit1:readdata -> mm_interconnect_0:digit1_s1_readdata
	wire   [2:0] mm_interconnect_0_digit1_s1_address;                          // mm_interconnect_0:digit1_s1_address -> digit1:address
	wire         mm_interconnect_0_digit1_s1_write;                            // mm_interconnect_0:digit1_s1_write -> digit1:write_n
	wire  [31:0] mm_interconnect_0_digit1_s1_writedata;                        // mm_interconnect_0:digit1_s1_writedata -> digit1:writedata
	wire         mm_interconnect_0_digit2_s1_chipselect;                       // mm_interconnect_0:digit2_s1_chipselect -> digit2:chipselect
	wire  [31:0] mm_interconnect_0_digit2_s1_readdata;                         // digit2:readdata -> mm_interconnect_0:digit2_s1_readdata
	wire   [2:0] mm_interconnect_0_digit2_s1_address;                          // mm_interconnect_0:digit2_s1_address -> digit2:address
	wire         mm_interconnect_0_digit2_s1_write;                            // mm_interconnect_0:digit2_s1_write -> digit2:write_n
	wire  [31:0] mm_interconnect_0_digit2_s1_writedata;                        // mm_interconnect_0:digit2_s1_writedata -> digit2:writedata
	wire         mm_interconnect_0_digit3_s1_chipselect;                       // mm_interconnect_0:digit3_s1_chipselect -> digit3:chipselect
	wire  [31:0] mm_interconnect_0_digit3_s1_readdata;                         // digit3:readdata -> mm_interconnect_0:digit3_s1_readdata
	wire   [2:0] mm_interconnect_0_digit3_s1_address;                          // mm_interconnect_0:digit3_s1_address -> digit3:address
	wire         mm_interconnect_0_digit3_s1_write;                            // mm_interconnect_0:digit3_s1_write -> digit3:write_n
	wire  [31:0] mm_interconnect_0_digit3_s1_writedata;                        // mm_interconnect_0:digit3_s1_writedata -> digit3:writedata
	wire         mm_interconnect_0_digit4_s1_chipselect;                       // mm_interconnect_0:digit4_s1_chipselect -> digit4:chipselect
	wire  [31:0] mm_interconnect_0_digit4_s1_readdata;                         // digit4:readdata -> mm_interconnect_0:digit4_s1_readdata
	wire   [2:0] mm_interconnect_0_digit4_s1_address;                          // mm_interconnect_0:digit4_s1_address -> digit4:address
	wire         mm_interconnect_0_digit4_s1_write;                            // mm_interconnect_0:digit4_s1_write -> digit4:write_n
	wire  [31:0] mm_interconnect_0_digit4_s1_writedata;                        // mm_interconnect_0:digit4_s1_writedata -> digit4:writedata
	wire         mm_interconnect_0_digit5_s1_chipselect;                       // mm_interconnect_0:digit5_s1_chipselect -> digit5:chipselect
	wire  [31:0] mm_interconnect_0_digit5_s1_readdata;                         // digit5:readdata -> mm_interconnect_0:digit5_s1_readdata
	wire   [2:0] mm_interconnect_0_digit5_s1_address;                          // mm_interconnect_0:digit5_s1_address -> digit5:address
	wire         mm_interconnect_0_digit5_s1_write;                            // mm_interconnect_0:digit5_s1_write -> digit5:write_n
	wire  [31:0] mm_interconnect_0_digit5_s1_writedata;                        // mm_interconnect_0:digit5_s1_writedata -> digit5:writedata
	wire         irq_mapper_receiver0_irq;                                     // opencores_i2c_0:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // pioPushButton:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                     // timer:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                         // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [digit0:reset_n, digit1:reset_n, digit2:reset_n, digit3:reset_n, digit4:reset_n, digit5:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory:reset, opencores_i2c_0:wb_rst_i, pioPushButton:reset_n, rst_translator:in_reset, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]

	lab3_qsys_digit0 digit0 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_digit0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_digit0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_digit0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_digit0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_digit0_s1_readdata),   //                    .readdata
		.out_port   (digit0_external_connection_export)       // external_connection.export
	);

	lab3_qsys_digit0 digit1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_digit1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_digit1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_digit1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_digit1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_digit1_s1_readdata),   //                    .readdata
		.out_port   (digit1_external_connection_export)       // external_connection.export
	);

	lab3_qsys_digit0 digit2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_digit2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_digit2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_digit2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_digit2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_digit2_s1_readdata),   //                    .readdata
		.out_port   (digit2_external_connection_export)       // external_connection.export
	);

	lab3_qsys_digit0 digit3 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_digit3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_digit3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_digit3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_digit3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_digit3_s1_readdata),   //                    .readdata
		.out_port   (digit3_external_connection_export)       // external_connection.export
	);

	lab3_qsys_digit0 digit4 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_digit4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_digit4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_digit4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_digit4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_digit4_s1_readdata),   //                    .readdata
		.out_port   (digit4_external_connection_export)       // external_connection.export
	);

	lab3_qsys_digit0 digit5 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_digit5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_digit5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_digit5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_digit5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_digit5_s1_readdata),   //                    .readdata
		.out_port   (digit5_external_connection_export)       // external_connection.export
	);

	lab3_qsys_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	lab3_qsys_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	lab3_qsys_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	opencores_i2c opencores_i2c_0 (
		.wb_clk_i   (clk_clk),                                                      //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                               //      clock_reset.reset
		.scl_pad_io (opencores_i2c_0_export_0_scl_pad_io),                          //         export_0.export
		.sda_pad_io (opencores_i2c_0_export_0_sda_pad_io),                          //                 .export
		.wb_adr_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                      // interrupt_sender.irq
	);

	lab3_qsys_pioPushButton piopushbutton (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_piopushbutton_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_piopushbutton_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_piopushbutton_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_piopushbutton_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_piopushbutton_s1_readdata),   //                    .readdata
		.in_port    (piopushbutton_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                       //                 irq.irq
	);

	lab3_qsys_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)               //   irq.irq
	);

	lab3_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                       //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                              //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                          //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                           //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                                 //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                             //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                                //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                            //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                          //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                       //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                   //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                          //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                      //                                         .readdata
		.digit0_s1_address                              (mm_interconnect_0_digit0_s1_address),                           //                                digit0_s1.address
		.digit0_s1_write                                (mm_interconnect_0_digit0_s1_write),                             //                                         .write
		.digit0_s1_readdata                             (mm_interconnect_0_digit0_s1_readdata),                          //                                         .readdata
		.digit0_s1_writedata                            (mm_interconnect_0_digit0_s1_writedata),                         //                                         .writedata
		.digit0_s1_chipselect                           (mm_interconnect_0_digit0_s1_chipselect),                        //                                         .chipselect
		.digit1_s1_address                              (mm_interconnect_0_digit1_s1_address),                           //                                digit1_s1.address
		.digit1_s1_write                                (mm_interconnect_0_digit1_s1_write),                             //                                         .write
		.digit1_s1_readdata                             (mm_interconnect_0_digit1_s1_readdata),                          //                                         .readdata
		.digit1_s1_writedata                            (mm_interconnect_0_digit1_s1_writedata),                         //                                         .writedata
		.digit1_s1_chipselect                           (mm_interconnect_0_digit1_s1_chipselect),                        //                                         .chipselect
		.digit2_s1_address                              (mm_interconnect_0_digit2_s1_address),                           //                                digit2_s1.address
		.digit2_s1_write                                (mm_interconnect_0_digit2_s1_write),                             //                                         .write
		.digit2_s1_readdata                             (mm_interconnect_0_digit2_s1_readdata),                          //                                         .readdata
		.digit2_s1_writedata                            (mm_interconnect_0_digit2_s1_writedata),                         //                                         .writedata
		.digit2_s1_chipselect                           (mm_interconnect_0_digit2_s1_chipselect),                        //                                         .chipselect
		.digit3_s1_address                              (mm_interconnect_0_digit3_s1_address),                           //                                digit3_s1.address
		.digit3_s1_write                                (mm_interconnect_0_digit3_s1_write),                             //                                         .write
		.digit3_s1_readdata                             (mm_interconnect_0_digit3_s1_readdata),                          //                                         .readdata
		.digit3_s1_writedata                            (mm_interconnect_0_digit3_s1_writedata),                         //                                         .writedata
		.digit3_s1_chipselect                           (mm_interconnect_0_digit3_s1_chipselect),                        //                                         .chipselect
		.digit4_s1_address                              (mm_interconnect_0_digit4_s1_address),                           //                                digit4_s1.address
		.digit4_s1_write                                (mm_interconnect_0_digit4_s1_write),                             //                                         .write
		.digit4_s1_readdata                             (mm_interconnect_0_digit4_s1_readdata),                          //                                         .readdata
		.digit4_s1_writedata                            (mm_interconnect_0_digit4_s1_writedata),                         //                                         .writedata
		.digit4_s1_chipselect                           (mm_interconnect_0_digit4_s1_chipselect),                        //                                         .chipselect
		.digit5_s1_address                              (mm_interconnect_0_digit5_s1_address),                           //                                digit5_s1.address
		.digit5_s1_write                                (mm_interconnect_0_digit5_s1_write),                             //                                         .write
		.digit5_s1_readdata                             (mm_interconnect_0_digit5_s1_readdata),                          //                                         .readdata
		.digit5_s1_writedata                            (mm_interconnect_0_digit5_s1_writedata),                         //                                         .writedata
		.digit5_s1_chipselect                           (mm_interconnect_0_digit5_s1_chipselect),                        //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),       //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),         //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),          //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),      //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),     //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),   //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),    //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),        //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),          //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),           //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),       //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),      //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),     //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),    //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),    //                                         .debugaccess
		.onchip_memory_s1_address                       (mm_interconnect_0_onchip_memory_s1_address),                    //                         onchip_memory_s1.address
		.onchip_memory_s1_write                         (mm_interconnect_0_onchip_memory_s1_write),                      //                                         .write
		.onchip_memory_s1_readdata                      (mm_interconnect_0_onchip_memory_s1_readdata),                   //                                         .readdata
		.onchip_memory_s1_writedata                     (mm_interconnect_0_onchip_memory_s1_writedata),                  //                                         .writedata
		.onchip_memory_s1_byteenable                    (mm_interconnect_0_onchip_memory_s1_byteenable),                 //                                         .byteenable
		.onchip_memory_s1_chipselect                    (mm_interconnect_0_onchip_memory_s1_chipselect),                 //                                         .chipselect
		.onchip_memory_s1_clken                         (mm_interconnect_0_onchip_memory_s1_clken),                      //                                         .clken
		.opencores_i2c_0_avalon_slave_0_address         (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_address),      //           opencores_i2c_0_avalon_slave_0.address
		.opencores_i2c_0_avalon_slave_0_write           (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_write),        //                                         .write
		.opencores_i2c_0_avalon_slave_0_readdata        (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_readdata),     //                                         .readdata
		.opencores_i2c_0_avalon_slave_0_writedata       (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_writedata),    //                                         .writedata
		.opencores_i2c_0_avalon_slave_0_waitrequest     (~mm_interconnect_0_opencores_i2c_0_avalon_slave_0_waitrequest), //                                         .waitrequest
		.opencores_i2c_0_avalon_slave_0_chipselect      (mm_interconnect_0_opencores_i2c_0_avalon_slave_0_chipselect),   //                                         .chipselect
		.pioPushButton_s1_address                       (mm_interconnect_0_piopushbutton_s1_address),                    //                         pioPushButton_s1.address
		.pioPushButton_s1_write                         (mm_interconnect_0_piopushbutton_s1_write),                      //                                         .write
		.pioPushButton_s1_readdata                      (mm_interconnect_0_piopushbutton_s1_readdata),                   //                                         .readdata
		.pioPushButton_s1_writedata                     (mm_interconnect_0_piopushbutton_s1_writedata),                  //                                         .writedata
		.pioPushButton_s1_chipselect                    (mm_interconnect_0_piopushbutton_s1_chipselect),                 //                                         .chipselect
		.timer_s1_address                               (mm_interconnect_0_timer_s1_address),                            //                                 timer_s1.address
		.timer_s1_write                                 (mm_interconnect_0_timer_s1_write),                              //                                         .write
		.timer_s1_readdata                              (mm_interconnect_0_timer_s1_readdata),                           //                                         .readdata
		.timer_s1_writedata                             (mm_interconnect_0_timer_s1_writedata),                          //                                         .writedata
		.timer_s1_chipselect                            (mm_interconnect_0_timer_s1_chipselect)                          //                                         .chipselect
	);

	lab3_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
